
`define PC_WIDTH            32
`define rv32_XLEN           32
`define RF_IDX_WIDTH        5
//`define RD_IDX_WIDTH        5
`define RF_REG_NUM          32
`define ADDIR0              `rv32_XLEN'h00000013

`define PC_add_insr         4
`define ADDRESS_rst         `PC_WIDTH'h00001000
`define address_sim         `ADDRESS_rst>>2

`define ADDR_Bpu_WIDTH      `PC_WIDTH     

    `define DECINFO_BJP_JUMP_LSB    0
    `define DECINFO_BJP_JUMP_MSB    `DECINFO_BJP_JUMP_LSB+1-1
`define DECINFO_BJP_JUMP            `DECINFO_BJP_JUMP_MSB:`DECINFO_BJP_JUMP_LSB
    `define DECINFO_BJP_BEQ_LSB     `DECINFO_BJP_JUMP_MSB+1
    `define DECINFO_BJP_BEQ_MSB     `DECINFO_BJP_BEQ_LSB+1-1
`define DECINFO_BJP_BEQ             `DECINFO_BJP_BEQ_MSB:`DECINFO_BJP_BEQ_LSB
    `define DECINFO_BJP_BNE_LSB     `DECINFO_BJP_BEQ_MSB+1
    `define DECINFO_BJP_BNE_MSB     `DECINFO_BJP_BNE_LSB+1-1
`define DECINFO_BJP_BNE             `DECINFO_BJP_BNE_MSB:`DECINFO_BJP_BNE_LSB
    `define DECINFO_BJP_BLT_LSB     `DECINFO_BJP_BNE_MSB+1
    `define DECINFO_BJP_BLT_MSB     `DECINFO_BJP_BLT_LSB+1-1
`define DECINFO_BJP_BLT             `DECINFO_BJP_BLT_MSB:`DECINFO_BJP_BLT_LSB
    `define DECINFO_BJP_BGT_LSB     `DECINFO_BJP_BLT_MSB+1
    `define DECINFO_BJP_BGT_MSB     `DECINFO_BJP_BGT_LSB+1-1
`define DECINFO_BJP_BGT             `DECINFO_BJP_BGT_MSB:`DECINFO_BJP_BGT_LSB
    `define DECINFO_BJP_BLTU_LSB    `DECINFO_BJP_BGT_MSB+1
    `define DECINFO_BJP_BLTU_MSB    `DECINFO_BJP_BLTU_LSB+1-1
`define DECINFO_BJP_BLTU            `DECINFO_BJP_BLTU_MSB:`DECINFO_BJP_BLTU_LSB
    `define DECINFO_BJP_BGTU_LSB    `DECINFO_BJP_BLTU_MSB+1
    `define DECINFO_BJP_BGTU_MSB    `DECINFO_BJP_BGTU_LSB+1-1
`define DECINFO_BJP_BGTU            `DECINFO_BJP_BGTU_MSB:`DECINFO_BJP_BGTU_LSB
    `define DECINFO_BJP_BXX_LSB     `DECINFO_BJP_BGTU_MSB+1
    `define DECINFO_BJP_BXX_MSB     `DECINFO_BJP_BXX_LSB+1-1
`define DECINFO_BJP_BXX             `DECINFO_BJP_BXX_MSB:`DECINFO_BJP_BXX_LSB
    `define DECINFO_BJP_FENCE_LSB   `DECINFO_BJP_BXX_MSB+1
    `define DECINFO_BJP_FENCE_MSB   `DECINFO_BJP_FENCE_LSB+1-1
`define DECINFO_BJP_FENCE           `DECINFO_BJP_FENCE_MSB:`DECINFO_BJP_FENCE_LSB
    `define DECINFO_BJP_FENCEI_LSB  `DECINFO_BJP_FENCE_MSB+1
    `define DECINFO_BJP_FENCEI_MSB  `DECINFO_BJP_FENCEI_LSB+1-1
`define DECINFO_BJP_FENCEI          `DECINFO_BJP_FENCEI_MSB:`DECINFO_BJP_FENCEI_LSB   
`define DECINFO_BJP_WIDTH           `DECINFO_BJP_FENCEI_MSB+1

    `define DECINFO_ALU_LSB         0
    `define DECINFO_ALU_MSB         `DECINFO_ALU_LSB+1-1
`define DECINFO_ALU                 `DECINFO_ALU_MSB:`DECINFO_ALU_LSB
    `define DECINFO_ALU_ADD_LSB     `DECINFO_ALU_MSB+1
    `define DECINFO_ALU_ADD_MSB     `DECINFO_ALU_ADD_LSB+1-1
`define DECINFO_ALU_ADD             `DECINFO_ALU_ADD_MSB:`DECINFO_ALU_ADD_LSB
    `define DECINFO_ALU_ADDI_LSB    `DECINFO_ALU_ADD_MSB+1
    `define DECINFO_ALU_ADDI_MSB    `DECINFO_ALU_ADDI_LSB+1-1
`define DECINFO_ALU_ADDI            `DECINFO_ALU_ADDI_MSB:`DECINFO_ALU_ADDI_LSB

    `define DECINFO_ALU_SUB_LSB     `DECINFO_ALU_ADDI_MSB+1
    `define DECINFO_ALU_SUB_MSB     `DECINFO_ALU_SUB_LSB+1-1
`define DECINFO_ALU_SUB             `DECINFO_ALU_SUB_MSB:`DECINFO_ALU_SUB_LSB
    `define DECINFO_ALU_SLT_LSB     `DECINFO_ALU_SUB_MSB+1
    `define DECINFO_ALU_SLT_MSB     `DECINFO_ALU_SLT_LSB+1-1
`define DECINFO_ALU_SLT             `DECINFO_ALU_SLT_MSB:`DECINFO_ALU_SLT_LSB
    `define DECINFO_ALU_SLTU_LSB    `DECINFO_ALU_SLT_MSB+1
    `define DECINFO_ALU_SLTU_MSB    `DECINFO_ALU_SLTU_LSB+1-1
`define DECINFO_ALU_SLTU            `DECINFO_ALU_SLTU_MSB:`DECINFO_ALU_SLTU_LSB
    `define DECINFO_ALU_SLTI_LSB    `DECINFO_ALU_SLTU_MSB+1
    `define DECINFO_ALU_SLTI_MSB    `DECINFO_ALU_SLTI_LSB+1-1
`define DECINFO_ALU_SLTI            `DECINFO_ALU_SLTI_MSB:`DECINFO_ALU_SLTI_LSB
    `define DECINFO_ALU_SLTIU_LSB   `DECINFO_ALU_SLTI_MSB+1
    `define DECINFO_ALU_SLTIU_MSB   `DECINFO_ALU_SLTIU_LSB+1-1
`define DECINFO_ALU_SLTIU           `DECINFO_ALU_SLTIU_MSB:`DECINFO_ALU_SLTIU_LSB
    `define DECINFO_ALU_XOR_LSB     `DECINFO_ALU_SLTIU_MSB+1
    `define DECINFO_ALU_XOR_MSB     `DECINFO_ALU_XOR_LSB+1-1
`define DECINFO_ALU_XOR             `DECINFO_ALU_XOR_MSB:`DECINFO_ALU_XOR_LSB
    `define DECINFO_ALU_XORI_LSB    `DECINFO_ALU_XOR_MSB+1
    `define DECINFO_ALU_XORI_MSB    `DECINFO_ALU_XORI_LSB+1-1
`define DECINFO_ALU_XORI            `DECINFO_ALU_XORI_MSB:`DECINFO_ALU_XORI_LSB

    `define DECINFO_ALU_SLL_LSB     `DECINFO_ALU_XORI_MSB+1
    `define DECINFO_ALU_SLL_MSB     `DECINFO_ALU_SLL_LSB+1-1
`define DECINFO_ALU_SLL             `DECINFO_ALU_SLL_MSB:`DECINFO_ALU_SLL_LSB
    `define DECINFO_ALU_SLLI_LSB    `DECINFO_ALU_SLL_MSB+1
    `define DECINFO_ALU_SLLI_MSB    `DECINFO_ALU_SLLI_LSB+1-1
`define DECINFO_ALU_SLLI            `DECINFO_ALU_SLLI_MSB:`DECINFO_ALU_SLLI_LSB

    `define DECINFO_ALU_SRL_LSB     `DECINFO_ALU_SLLI_MSB+1
    `define DECINFO_ALU_SRL_MSB     `DECINFO_ALU_SRL_LSB+1-1
`define DECINFO_ALU_SRL             `DECINFO_ALU_SRL_MSB:`DECINFO_ALU_SRL_LSB
    `define DECINFO_ALU_SRLI_LSB    `DECINFO_ALU_SRL_MSB+1
    `define DECINFO_ALU_SRLI_MSB    `DECINFO_ALU_SRLI_LSB+1-1
`define DECINFO_ALU_SRLI            `DECINFO_ALU_SRLI_MSB:`DECINFO_ALU_SRLI_LSB


    `define DECINFO_ALU_SRA_LSB     `DECINFO_ALU_SRLI_MSB+1
    `define DECINFO_ALU_SRA_MSB     `DECINFO_ALU_SRA_LSB+1-1
`define DECINFO_ALU_SRA             `DECINFO_ALU_SRA_MSB:`DECINFO_ALU_SRA_LSB
    `define DECINFO_ALU_SRAI_LSB    `DECINFO_ALU_SRA_MSB+1
    `define DECINFO_ALU_SRAI_MSB    `DECINFO_ALU_SRAI_LSB+1-1
`define DECINFO_ALU_SRAI            `DECINFO_ALU_SRAI_MSB:`DECINFO_ALU_SRAI_LSB

    `define DECINFO_ALU_OR_LSB      `DECINFO_ALU_SRAI_MSB+1
    `define DECINFO_ALU_OR_MSB      `DECINFO_ALU_OR_LSB+1-1
`define DECINFO_ALU_OR              `DECINFO_ALU_OR_MSB:`DECINFO_ALU_OR_LSB
    `define DECINFO_ALU_ORI_LSB     `DECINFO_ALU_OR_MSB+1
    `define DECINFO_ALU_ORI_MSB     `DECINFO_ALU_ORI_LSB+1-1
`define DECINFO_ALU_ORI             `DECINFO_ALU_ORI_MSB:`DECINFO_ALU_ORI_LSB


    `define DECINFO_ALU_AND_LSB     `DECINFO_ALU_ORI_MSB+1
    `define DECINFO_ALU_AND_MSB     `DECINFO_ALU_AND_LSB+1-1
`define DECINFO_ALU_AND             `DECINFO_ALU_AND_MSB:`DECINFO_ALU_AND_LSB
    `define DECINFO_ALU_ANDI_LSB    `DECINFO_ALU_AND_MSB+1
    `define DECINFO_ALU_ANDI_MSB    `DECINFO_ALU_ANDI_LSB+1-1
`define DECINFO_ALU_ANDI            `DECINFO_ALU_ANDI_MSB:`DECINFO_ALU_ANDI_LSB

    `define DECINFO_ALU_LUI_LSB     `DECINFO_ALU_ANDI_MSB+1
    `define DECINFO_ALU_LUI_MSB     `DECINFO_ALU_LUI_LSB+1-1
`define DECINFO_ALU_LUI             `DECINFO_ALU_LUI_MSB:`DECINFO_ALU_LUI_LSB
    `define DECINFO_ALU_auipc_LSB   `DECINFO_ALU_LUI_MSB+1
    `define DECINFO_ALU_auipc_MSB   `DECINFO_ALU_auipc_LSB+1-1
`define DECINFO_ALU_auipc           `DECINFO_ALU_auipc_MSB:`DECINFO_ALU_auipc_LSB
    `define DECINFO_ALU_NOP_LSB     `DECINFO_ALU_auipc_MSB+1
    `define DECINFO_ALU_NOP_MSB     `DECINFO_ALU_NOP_LSB+1-1
`define DECINFO_ALU_NOP             `DECINFO_ALU_NOP_MSB:`DECINFO_ALU_NOP_LSB
    `define DECINFO_ALU_ECAL_LSB    `DECINFO_ALU_NOP_MSB+1
    `define DECINFO_ALU_ECAL_MSB    `DECINFO_ALU_ECAL_LSB+1-1
`define DECINFO_ALU_ECAL            `DECINFO_ALU_ECAL_MSB:`DECINFO_ALU_ECAL_LSB
    `define DECINFO_ALU_EBRK_LSB    `DECINFO_ALU_ECAL_MSB+1
    `define DECINFO_ALU_EBRK_MSB    `DECINFO_ALU_EBRK_LSB+1-1
`define DECINFO_ALU_EBRK            `DECINFO_ALU_EBRK_MSB:`DECINFO_ALU_EBRK_LSB
`define DECINFO_ALU_WIDTH           `DECINFO_ALU_EBRK_MSB+1


`define DECINFO_CSR_CSRRW           0   
`define DECINFO_CSR_CSRRS           `DECINFO_CSR_CSRRW+1
`define DECINFO_CSR_CSRRC           `DECINFO_CSR_CSRRS+1
`define DECINFO_CSR_WIDTH           `DECINFO_CSR_CSRRC+1

    `define DECINFO_L_S_LSB         0
    `define DECINFO_L_S_MSB         `DECINFO_L_S_LSB+1-1
`define DECINFO_L_S                 `DECINFO_L_S_MSB:`DECINFO_L_S_LSB
    `define DECINFO_LOAD_LB_LSB     `DECINFO_L_S_MSB+1
    `define DECINFO_LOAD_LB_MSB     `DECINFO_LOAD_LB_LSB+1-1
`define DECINFO_LOAD_LB             `DECINFO_LOAD_LB_MSB:`DECINFO_LOAD_LB_LSB
    `define DECINFO_LOAD_LH_LSB     `DECINFO_LOAD_LB_MSB+1
    `define DECINFO_LOAD_LH_MSB     `DECINFO_LOAD_LH_LSB+1-1
`define DECINFO_LOAD_LH             `DECINFO_LOAD_LH_MSB:`DECINFO_LOAD_LH_LSB
    `define DECINFO_LOAD_LW_LSB     `DECINFO_LOAD_LH_MSB+1
    `define DECINFO_LOAD_LW_MSB     `DECINFO_LOAD_LW_LSB+1-1
`define DECINFO_LOAD_LW             `DECINFO_LOAD_LW_MSB:`DECINFO_LOAD_LW_LSB
    `define DECINFO_LOAD_LBU_LSB    `DECINFO_LOAD_LW_MSB+1
    `define DECINFO_LOAD_LBU_MSB    `DECINFO_LOAD_LBU_LSB+1-1
`define DECINFO_LOAD_LBU            `DECINFO_LOAD_LBU_MSB:`DECINFO_LOAD_LBU_LSB
    `define DECINFO_LOAD_LHU_LSB    `DECINFO_LOAD_LBU_MSB+1
    `define DECINFO_LOAD_LHU_MSB    `DECINFO_LOAD_LHU_LSB+1-1
`define DECINFO_LOAD_LHU            `DECINFO_LOAD_LHU_MSB:`DECINFO_LOAD_LHU_LSB
    `define DECINFO_Stor_SB_LSB     `DECINFO_LOAD_LHU_MSB+1
    `define DECINFO_Stor_SB_MSB     `DECINFO_Stor_SB_LSB+1-1
`define DECINFO_Stor_SB             `DECINFO_Stor_SB_MSB:`DECINFO_Stor_SB_LSB
    `define DECINFO_Stor_SH_LSB     `DECINFO_Stor_SB_MSB+1
    `define DECINFO_Stor_SH_MSB     `DECINFO_Stor_SH_LSB+1-1
`define DECINFO_Stor_SH             `DECINFO_Stor_SH_MSB:`DECINFO_Stor_SH_LSB
    `define DECINFO_Stor_SW_LSB     `DECINFO_Stor_SH_MSB+1
    `define DECINFO_Stor_SW_MSB     `DECINFO_Stor_SW_LSB+1-1
`define DECINFO_Stor_SW             `DECINFO_Stor_SW_MSB:`DECINFO_Stor_SW_LSB
`define DECINFO_L_S_WIDTH           `DECINFO_Stor_SW_MSB+1
   
    `define DECINFO_MD_LSB          0
    `define DECINFO_MD_MSB          `DECINFO_MD_LSB+1-1
`define DECINFO_MD                  `DECINFO_MD_MSB:`DECINFO_MD_LSB
    `define DECINFO_MD_MUL_LSB      `DECINFO_MD_MSB+1
    `define DECINFO_MD_MUL_MSB      `DECINFO_MD_MUL_LSB+1-1
`define DECINFO_MD_MUL              `DECINFO_MD_MUL_MSB:`DECINFO_MD_MUL_LSB
    `define DECINFO_MD_MULH_LSB     `DECINFO_MD_MUL_MSB+1
    `define DECINFO_MD_MULH_MSB     `DECINFO_MD_MULH_LSB+1-1
`define DECINFO_MD_MULH             `DECINFO_MD_MULH_MSB:`DECINFO_MD_MULH_LSB
    `define DECINFO_MD_MULHU_LSB    `DECINFO_MD_MULH_MSB+1
    `define DECINFO_MD_MULHU_MSB    `DECINFO_MD_MULHU_LSB+1-1
`define DECINFO_MD_MULHU            `DECINFO_MD_MULHU_MSB:`DECINFO_MD_MULHU_LSB
    `define DECINFO_MD_MULHSU_LSB   `DECINFO_MD_MULHU_MSB+1
    `define DECINFO_MD_MULHSU_MSB   `DECINFO_MD_MULHSU_LSB+1-1
`define DECINFO_MD_MULHSU           `DECINFO_MD_MULHSU_MSB:`DECINFO_MD_MULHSU_LSB
    `define DECINFO_MUL_LSB         `DECINFO_MD_MULHSU_MSB+1
    `define DECINFO_MUL_MSB         `DECINFO_MUL_LSB+1-1
`define DECINFO_MUL                 `DECINFO_MUL_MSB:`DECINFO_MUL_LSB
    `define DECINFO_MD_DIV_LSB      `DECINFO_MUL_MSB+1
    `define DECINFO_MD_DIV_MSB      `DECINFO_MD_DIV_LSB+1-1
`define DECINFO_MD_DIV              `DECINFO_MD_DIV_MSB:`DECINFO_MD_DIV_LSB
    `define DECINFO_MD_DIVU_LSB     `DECINFO_MD_DIV_MSB+1
    `define DECINFO_MD_DIVU_MSB     `DECINFO_MD_DIVU_LSB+1-1
`define DECINFO_MD_DIVU             `DECINFO_MD_DIVU_MSB:`DECINFO_MD_DIVU_LSB
    `define DECINFO_MD_REM_LSB      `DECINFO_MD_DIVU_MSB+1
    `define DECINFO_MD_REM_MSB      `DECINFO_MD_REM_LSB+1-1
`define DECINFO_MD_REM              `DECINFO_MD_REM_MSB:`DECINFO_MD_REM_LSB
    `define DECINFO_MD_REMU_LSB     `DECINFO_MD_REM_MSB+1
    `define DECINFO_MD_REMU_MSB     `DECINFO_MD_REMU_LSB+1-1
`define DECINFO_MD_REMU             `DECINFO_MD_REMU_MSB:`DECINFO_MD_REMU_LSB
    `define DECINFO_DIV_LSB         `DECINFO_MD_REMU_MSB+1
    `define DECINFO_DIV_MSB         `DECINFO_DIV_LSB+1-1
`define DECINFO_DIV                 `DECINFO_DIV_MSB:`DECINFO_DIV_LSB
`define DECINFO_M_D_WIDTH           `DECINFO_DIV_MSB+1

    `define add_en                  0
    `define com_en                  `add_en+1
    `define and_en                  `com_en+1
    `define or_en                   `and_en+1
    `define xor_en                  `or_en+1
    `define lgcl_en                 `xor_en+1
    `define lgc_en                  `lgcl_en+1
    `define alur_en                 `lgc_en+1
    //`define mul_en                  `alur_en+1
    //`define div_en                  `mul_en+1
    `define com_sign                `alur_en+1
    //`define lui_en                  `div_en+1
    `define EN_Wid                  `com_sign+1